module _4zm16decoder (clk, rst, Ind, En, \4 , \5 , \6 , \7 , \0 , \1 , \2 , \3 , \8 , \9 , \10 , \11 , \15 , \14 , \13 , \12 );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Ind;
  input  wire [0:0] En;
  output  wire [0:0] \4 ;
  output  wire [0:0] \5 ;
  output  wire [0:0] \6 ;
  output  wire [0:0] \7 ;
  output  wire [0:0] \0 ;
  output  wire [0:0] \1 ;
  output  wire [0:0] \2 ;
  output  wire [0:0] \3 ;
  output  wire [0:0] \8 ;
  output  wire [0:0] \9 ;
  output  wire [0:0] \10 ;
  output  wire [0:0] \11 ;
  output  wire [0:0] \15 ;
  output  wire [0:0] \14 ;
  output  wire [0:0] \13 ;
  output  wire [0:0] \12 ;

  TC_Splitter8 # (.UUID(64'd2846459251964735202 ^ UUID)) Splitter8_0 (.in(wire_3), .out0(wire_14), .out1(wire_1), .out2(wire_4), .out3(wire_5), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd445380417365926464 ^ UUID)) Decoder3_1 (.dis(wire_10), .sel0(wire_14), .sel1(wire_1), .sel2(wire_4), .out0(wire_18), .out1(wire_9), .out2(wire_23), .out3(wire_17), .out4(wire_22), .out5(wire_7), .out6(wire_28), .out7(wire_26));
  TC_Splitter8 # (.UUID(64'd4132815552358996771 ^ UUID)) Splitter8_2 (.in(wire_3), .out0(wire_27), .out1(wire_13), .out2(wire_12), .out3(wire_25), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd4403838804956136719 ^ UUID)) Decoder3_3 (.dis(wire_21), .sel0(wire_27), .sel1(wire_13), .sel2(wire_12), .out0(wire_29), .out1(wire_8), .out2(wire_16), .out3(wire_20), .out4(wire_0), .out5(wire_11), .out6(wire_19), .out7(wire_2));
  TC_Not # (.UUID(64'd4179574134841425537 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_25), .out(wire_6));
  TC_Not # (.UUID(64'd1850851141294105609 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_15), .out(wire_24));
  TC_Or # (.UUID(64'd464008523248432561 ^ UUID), .BIT_WIDTH(64'd1)) Or_6 (.in0(wire_24), .in1(wire_5), .out(wire_10));
  TC_Or # (.UUID(64'd2604936541790780610 ^ UUID), .BIT_WIDTH(64'd1)) Or_7 (.in0(wire_6), .in1(wire_24), .out(wire_21));
  TC_Constant # (.UUID(64'd1817809215004476502 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_8 (.out());
  TC_Constant # (.UUID(64'd4500563200943663130 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_9 (.out());
  TC_Constant # (.UUID(64'd4553730726826982281 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_10 (.out());
  TC_Constant # (.UUID(64'd2676911755365734023 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_11 (.out());
  TC_Constant # (.UUID(64'd2293009349816174489 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_12 (.out());
  TC_Constant # (.UUID(64'd4150386907538013779 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_13 (.out());
  TC_Constant # (.UUID(64'd1052125708879918401 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_14 (.out());
  TC_Constant # (.UUID(64'd287476249922060092 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_15 (.out());

  wire [0:0] wire_0;
  assign \12  = wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign \15  = wire_2;
  wire [7:0] wire_3;
  assign wire_3 = Ind;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign \5  = wire_7;
  wire [0:0] wire_8;
  assign \9  = wire_8;
  wire [0:0] wire_9;
  assign \1  = wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  assign \13  = wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  assign wire_15 = En;
  wire [0:0] wire_16;
  assign \10  = wire_16;
  wire [0:0] wire_17;
  assign \3  = wire_17;
  wire [0:0] wire_18;
  assign \0  = wire_18;
  wire [0:0] wire_19;
  assign \14  = wire_19;
  wire [0:0] wire_20;
  assign \11  = wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  assign \4  = wire_22;
  wire [0:0] wire_23;
  assign \2  = wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  assign \7  = wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  assign \6  = wire_28;
  wire [0:0] wire_29;
  assign \8  = wire_29;

endmodule
