module RegisterGroup (clk, rst, In_addr, Out_addr1, Out_addr2, En_In, Data_in, Out1_sbit7, Out1_sbit6, In_sbit6, In_sbit7, Out2_sbit6, Out2_sbit7, Data_out1, Data_out2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] In_addr;
  input  wire [7:0] Out_addr1;
  input  wire [7:0] Out_addr2;
  input  wire [0:0] En_In;
  input  wire [7:0] Data_in;
  output  wire [0:0] Out1_sbit7;
  output  wire [0:0] Out1_sbit6;
  output  wire [0:0] In_sbit6;
  output  wire [0:0] In_sbit7;
  output  wire [0:0] Out2_sbit6;
  output  wire [0:0] Out2_sbit7;
  output  wire [7:0] Data_out1;
  output  wire [7:0] Data_out2;

  TC_Constant # (.UUID(64'd2476018436133498686 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_0 (.out());
  TC_Constant # (.UUID(64'd2168569963486479072 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_1 (.out());
  TC_Constant # (.UUID(64'd4043736217543807666 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_2 (.out());
  TC_Constant # (.UUID(64'd396542217003720953 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_3 (.out());
  TC_Constant # (.UUID(64'd3954867635762248856 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_4 (.out());
  TC_Nor # (.UUID(64'd2084898473450824506 ^ UUID), .BIT_WIDTH(64'd1)) Nor_5 (.in0(wire_10), .in1(wire_17), .out(wire_24));
  TC_Nor # (.UUID(64'd1141109289603326753 ^ UUID), .BIT_WIDTH(64'd1)) Nor_6 (.in0(wire_43), .in1(wire_22), .out(wire_53));
  TC_Switch # (.UUID(64'd525243077953246989 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_36), .in(wire_56), .out(wire_4));
  TC_Nor # (.UUID(64'd2914653035550825021 ^ UUID), .BIT_WIDTH(64'd1)) Nor_8 (.in0(wire_7), .in1(wire_12), .out(wire_36));
  TC_Switch # (.UUID(64'd4529065468593763085 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_9 (.en(wire_53), .in(wire_1), .out(Data_out1));
  TC_Switch # (.UUID(64'd4138164610443691443 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_10 (.en(wire_24), .in(wire_0), .out(Data_out2));
  TC_Constant # (.UUID(64'd2317704081270560087 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_11 (.out());
  TC_Constant # (.UUID(64'd1316617174038851627 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_12 (.out());
  TC_Constant # (.UUID(64'd2780613661773122766 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_50));
  TC_Constant # (.UUID(64'd383966840177983124 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_57));
  _4zm16decoder # (.UUID(64'd1523080043891880085 ^ UUID)) _4zm16decoder_15 (.clk(clk), .rst(rst), .Ind(wire_46), .En(wire_9), .\4 (wire_48), .\5 (wire_2), .\6 (wire_7), .\7 (wire_12), .\0 (wire_13), .\1 (wire_6), .\2 (wire_52), .\3 (wire_40), .\8 (wire_14), .\9 (wire_21), .\10 (wire_60), .\11 (wire_19), .\15 (wire_20), .\14 (wire_35), .\13 (wire_45), .\12 (wire_49));
  _4zm16decoder # (.UUID(64'd3465023552995234528 ^ UUID)) _4zm16decoder_16 (.clk(clk), .rst(rst), .Ind(wire_16), .En(wire_57), .\4 (wire_38), .\5 (wire_31), .\6 (wire_43), .\7 (wire_22), .\0 (wire_23), .\1 (wire_39), .\2 (wire_25), .\3 (wire_29), .\8 (wire_41), .\9 (wire_8), .\10 (wire_15), .\11 (wire_32), .\15 (wire_3), .\14 (wire_18), .\13 (wire_26), .\12 (wire_5));
  RegisterPro # (.UUID(64'd3486757274636192172 ^ UUID)) RegisterPro_17 (.clk(clk), .rst(rst), .s1(wire_29), .s2(wire_42), .\�___________ (wire_4), .\�_____ (wire_40), .Out1(wire_1_5), .Out2(wire_0_8));
  RegisterPro # (.UUID(64'd4148574735080963847 ^ UUID)) RegisterPro_18 (.clk(clk), .rst(rst), .s1(wire_25), .s2(wire_55), .\�___________ (wire_4), .\�_____ (wire_52), .Out1(wire_1_8), .Out2(wire_0_10));
  RegisterPro # (.UUID(64'd1805533346382495819 ^ UUID)) RegisterPro_19 (.clk(clk), .rst(rst), .s1(wire_39), .s2(wire_33), .\�___________ (wire_4), .\�_____ (wire_6), .Out1(wire_1_13), .Out2(wire_0_12));
  RegisterPro # (.UUID(64'd1226882864486211718 ^ UUID)) RegisterPro_20 (.clk(clk), .rst(rst), .s1(wire_23), .s2(wire_44), .\�___________ (wire_4), .\�_____ (wire_13), .Out1(wire_1_12), .Out2(wire_0_13));
  RegisterPro # (.UUID(64'd1564765681901882392 ^ UUID)) RegisterPro_21 (.clk(clk), .rst(rst), .s1(wire_38), .s2(wire_27), .\�___________ (wire_4), .\�_____ (wire_48), .Out1(wire_1_14), .Out2(wire_0_14));
  RegisterPro # (.UUID(64'd4343002892340607771 ^ UUID)) RegisterPro_22 (.clk(clk), .rst(rst), .s1(wire_31), .s2(wire_54), .\�___________ (wire_4), .\�_____ (wire_2), .Out1(wire_1_15), .Out2(wire_0_15));
  RegisterPro # (.UUID(64'd3139442232711950001 ^ UUID)) RegisterPro_23 (.clk(clk), .rst(rst), .s1(wire_41), .s2(wire_30), .\�___________ (wire_4), .\�_____ (wire_14), .Out1(wire_1_9), .Out2(wire_0_11));
  RegisterPro # (.UUID(64'd330839372662474781 ^ UUID)) RegisterPro_24 (.clk(clk), .rst(rst), .s1(wire_8), .s2(wire_59), .\�___________ (wire_4), .\�_____ (wire_21), .Out1(wire_1_6), .Out2(wire_0_9));
  RegisterPro # (.UUID(64'd2893214525367273806 ^ UUID)) RegisterPro_25 (.clk(clk), .rst(rst), .s1(wire_26), .s2(wire_34), .\�___________ (wire_4), .\�_____ (wire_45), .Out1(wire_1_4), .Out2(wire_0_4));
  RegisterPro # (.UUID(64'd3368357102663641886 ^ UUID)) RegisterPro_26 (.clk(clk), .rst(rst), .s1(wire_5), .s2(wire_28), .\�___________ (wire_4), .\�_____ (wire_49), .Out1(wire_1_7), .Out2(wire_0_3));
  RegisterPro # (.UUID(64'd1747880564949271934 ^ UUID)) RegisterPro_27 (.clk(clk), .rst(rst), .s1(wire_32), .s2(wire_37), .\�___________ (wire_4), .\�_____ (wire_19), .Out1(wire_1_10), .Out2(wire_0_0));
  RegisterPro # (.UUID(64'd2632434431032018289 ^ UUID)) RegisterPro_28 (.clk(clk), .rst(rst), .s1(wire_15), .s2(wire_58), .\�___________ (wire_4), .\�_____ (wire_60), .Out1(wire_1_11), .Out2(wire_0_2));
  RegisterPro # (.UUID(64'd1608385328113584633 ^ UUID)) RegisterPro_29 (.clk(clk), .rst(rst), .s1(wire_18), .s2(wire_51), .\�___________ (wire_4), .\�_____ (wire_35), .Out1(wire_1_3), .Out2(wire_0_1));
  RegisterPro # (.UUID(64'd3453607857538586617 ^ UUID)) RegisterPro_30 (.clk(clk), .rst(rst), .s1(wire_3), .s2(wire_47), .\�___________ (wire_4), .\�_____ (wire_20), .Out1(wire_1_2), .Out2(wire_0_6));
  RegisterPro # (.UUID(64'd3303532811907655170 ^ UUID)) RegisterPro_31 (.clk(clk), .rst(rst), .s1(1'd0), .s2(1'd0), .\�___________ (wire_4), .\�_____ (1'd0), .Out1(wire_1_0), .Out2(wire_0_5));
  RegisterPro # (.UUID(64'd2001900293685094634 ^ UUID)) RegisterPro_32 (.clk(clk), .rst(rst), .s1(1'd0), .s2(1'd0), .\�___________ (wire_4), .\�_____ (1'd0), .Out1(wire_1_1), .Out2(wire_0_7));
  _4zm16decoder # (.UUID(64'd3244369760561604386 ^ UUID)) _4zm16decoder_33 (.clk(clk), .rst(rst), .Ind(wire_11), .En(wire_50), .\4 (wire_27), .\5 (wire_54), .\6 (wire_17), .\7 (wire_10), .\0 (wire_44), .\1 (wire_33), .\2 (wire_55), .\3 (wire_42), .\8 (wire_30), .\9 (wire_59), .\10 (wire_58), .\11 (wire_37), .\15 (wire_47), .\14 (wire_51), .\13 (wire_34), .\12 (wire_28));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  wire [7:0] wire_0_4;
  wire [7:0] wire_0_5;
  wire [7:0] wire_0_6;
  wire [7:0] wire_0_7;
  wire [7:0] wire_0_8;
  wire [7:0] wire_0_9;
  wire [7:0] wire_0_10;
  wire [7:0] wire_0_11;
  wire [7:0] wire_0_12;
  wire [7:0] wire_0_13;
  wire [7:0] wire_0_14;
  wire [7:0] wire_0_15;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6|wire_0_7|wire_0_8|wire_0_9|wire_0_10|wire_0_11|wire_0_12|wire_0_13|wire_0_14|wire_0_15;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  wire [7:0] wire_1_2;
  wire [7:0] wire_1_3;
  wire [7:0] wire_1_4;
  wire [7:0] wire_1_5;
  wire [7:0] wire_1_6;
  wire [7:0] wire_1_7;
  wire [7:0] wire_1_8;
  wire [7:0] wire_1_9;
  wire [7:0] wire_1_10;
  wire [7:0] wire_1_11;
  wire [7:0] wire_1_12;
  wire [7:0] wire_1_13;
  wire [7:0] wire_1_14;
  wire [7:0] wire_1_15;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8|wire_1_9|wire_1_10|wire_1_11|wire_1_12|wire_1_13|wire_1_14|wire_1_15;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign In_sbit6 = wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  assign wire_9 = En_In;
  wire [0:0] wire_10;
  assign Out2_sbit7 = wire_10;
  wire [7:0] wire_11;
  assign wire_11 = Out_addr2;
  wire [0:0] wire_12;
  assign In_sbit7 = wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  assign wire_16 = Out_addr1;
  wire [0:0] wire_17;
  assign Out2_sbit6 = wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  assign Out1_sbit7 = wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  assign Out1_sbit6 = wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [7:0] wire_46;
  assign wire_46 = In_addr;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  assign wire_56 = Data_in;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;

endmodule
